module multiplier(input logic Clk, Reset, Run, ClearA_LoadB,
					output [7:0]  Aval,    		
                                Bval,    		
                  output [6:0]  AhexL,			
                                AhexU,
                                BhexU,
                                BhexL,
                   output logic X
);





endmodule