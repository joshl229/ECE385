module processor(input logic	clk,
										[7:0] s, 
										reset, 
										run,
										cleara_loadb,
						
						output logic [6:0] ahexu, ahexl, bhexu, bhexl,
						output logic [7:0] aval, bval,
						output logic x);
						
// 						
						
										
										
							